module bitty(
    
);
endmodule;