/*
1111
0111
0011
*/